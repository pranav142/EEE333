module ALU_tb();
endmodule


