module error(input A, output F); 
assign A = 1'b0;
assign A = 1'b1;
assign F = A;
endmodule
