// 1. FIGURE OUT WHAT THE PROGRAM DOES!!!

module reg_file();

endmodule
